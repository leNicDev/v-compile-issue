module main

import calculator

fn main() {
        result := calculator,add(1, 2)
	println('1 + 2 = ${result}')
}
