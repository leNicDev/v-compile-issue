module calculator

pub fn add(a int, b int) {
  return a + b
}
